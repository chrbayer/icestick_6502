// tst_6502.v - test 6502 core
// 02-11-19 E. Brombaugh

module soc_6502(
    input clk,              // 4..0MHz CPU clock
    input reset,            // Low-true reset

	output reg [7:0] gpio_o,
	input [7:0] gpio_i,

	input RX,				// serial RX
	output TX				// serial TX
);
    // The 6502
    wire [15:0] CPU_AB;
    reg [7:0] CPU_DI;
    wire [7:0] CPU_DO;
    wire CPU_WE, CPU_IRQ;
    cpu_65ce02 ucpu(
        .clk(clk),
        .reset(reset),
        .AB(CPU_AB),
        .DI(CPU_DI),
        .DO(CPU_DO),
        .WE(CPU_WE),
        .IRQ(CPU_IRQ),
        .NMI(1'b0),
        .RDY(1'b1)
    );

	// address decode - not fully decoded for 512-byte memories
	wire p0 = (CPU_AB[15:12] == 4'h0) ? 1 : 0;
	wire p1 = (CPU_AB[15:12] == 4'h1) ? 1 : 0;
	wire p2 = (CPU_AB[15:12] == 4'h2) ? 1 : 0;
	wire pf = (CPU_AB[15:12] == 4'hf) ? 1 : 0;

	// RAM @ pages 00-0f
	reg [7:0] ram_mem [0:4095];
	initial
        $readmemh("null.hex", ram_mem);
	reg [7:0] ram_do;
	always @(posedge clk)
		if((CPU_WE == 1'b1) && (p0 == 1'b1))
			ram_mem[CPU_AB[11:0]] <= CPU_DO;
	always @(posedge clk)
		ram_do <= ram_mem[CPU_AB[11:0]];

	// CIA @ page 10-1f
	reg phi2;
	reg [7:0] cia_do;
	reg irq_n;
	reg [7:0] pa_out;
	reg [7:0] pb_in;
	reg flag_n;
	reg pc_n;
	reg tod;
	reg sp_in;
	reg sp_out;
	reg cnt_in;
	reg cnt_out;
	mos6526 umos6526(
		.clk(clk),
		.phi2(phi2), // Phi 2 positive edge
		.res_n(~reset),
		.cs_n(~p1),
		.rw(CPU_WE),
		.rs(CPU_AB[3:0]),
		.db_in(CPU_DO),
		.db_out(cia_do),
		.pa_in(gpio_i),
		.pa_out(pa_out),
		.pb_in(pb_in),
		.pb_out(gpio_o),
		.flag_n(flag_n),
		.pc_n(pc_n),
		.tod(tod),
		.sp_in(sp_in),
		.sp_out(sp_out),
		.cnt_in(cnt_in),
		.cnt_out(cnt_out),
		.irq_n(irq_n)
	);

	// ACIA at page 20-2f
	wire [7:0] acia_do;
	acia uacia(
		.clk(clk),				// system clock
		.rst(reset),			// system reset
		.cs(p2),				// chip select
		.we(CPU_WE),			// write enable
		.rs(CPU_AB[0]),			// register select
		.rx(RX),				// serial receive
		.din(CPU_DO),			// data bus input
		.dout(acia_do),			// data bus output
		.tx(TX),				// serial transmit
		.irq(CPU_IRQ)			// interrupt request
	);

	// ROM @ pages f0,f1...
	reg [7:0] rom_do;
`ifdef VERIFICATION
    reg [7:0] rom_mem [0:16383];
	initial
`ifdef VERIFICATION_6502
        $readmemh("6502_verification.hex", rom_mem);
`endif
`ifdef VERIFICATION_65C02
        $readmemh("65C02_verification.hex", rom_mem);
`endif
`ifdef DECIMAL_TEST_65C02
        $readmemh("65C02_decimal_test.hex", rom_mem);
`endif
`ifdef VERIFICATION_65CE02
        $readmemh("65CE02_opcodes_test.hex", rom_mem);
`endif
	always @(posedge clk)
		rom_do <= rom_mem[CPU_AB[13:0]];
`ifdef SIM
	initial
`ifdef VERIFICATION_6502
		$monitor("#%0t test_case = %0h", $time, ram_mem[512]);
`endif
`ifdef VERIFICATION_65C02
		$monitor("#%0t test_case = %0h", $time, ram_mem[512]);
`endif
`ifdef DECIMAL_TEST_65C02
		$monitor("#%0t ERROR = %0h", $time, ram_mem[11]);
`endif
`ifdef VERIFICATION_65CE02
		$monitor("#%0t test_case = %0h", $time, ram_mem[514]);
`endif
`endif
`else
    reg [7:0] rom_mem [0:4095];
	initial
        $readmemh("rom.hex", rom_mem);
	always @(posedge clk)
		rom_do <= rom_mem[CPU_AB[11:0]];
`endif


	// data mux
	reg [3:0] mux_sel;
	always @(posedge clk)
		mux_sel <= CPU_AB[15:12];
	always @(*)
		casez(mux_sel)
			4'h0: CPU_DI = ram_do;
			4'h1: CPU_DI = cia_do;
			4'h2: CPU_DI = acia_do;
			4'hf: CPU_DI = rom_do;
			default: CPU_DI = rom_do;
		endcase
endmodule
